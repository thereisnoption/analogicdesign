magic
tech sky130A
magscale 1 2
timestamp 1729238048
<< nmos >>
rect -189 -100 -29 100
rect 29 -100 189 100
<< ndiff >>
rect -247 88 -189 100
rect -247 -88 -235 88
rect -201 -88 -189 88
rect -247 -100 -189 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 189 88 247 100
rect 189 -88 201 88
rect 235 -88 247 88
rect 189 -100 247 -88
<< ndiffc >>
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
<< poly >>
rect -189 172 -29 188
rect -189 138 -173 172
rect -45 138 -29 172
rect -189 100 -29 138
rect 29 172 189 188
rect 29 138 45 172
rect 173 138 189 172
rect 29 100 189 138
rect -189 -138 -29 -100
rect -189 -172 -173 -138
rect -45 -172 -29 -138
rect -189 -188 -29 -172
rect 29 -138 189 -100
rect 29 -172 45 -138
rect 173 -172 189 -138
rect 29 -188 189 -172
<< polycont >>
rect -173 138 -45 172
rect 45 138 173 172
rect -173 -172 -45 -138
rect 45 -172 173 -138
<< locali >>
rect -189 138 -173 172
rect -45 138 -29 172
rect 29 138 45 172
rect 173 138 189 172
rect -235 88 -201 104
rect -235 -104 -201 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 201 88 235 104
rect 201 -104 235 -88
rect -189 -172 -173 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 173 -172 189 -138
<< viali >>
rect -160 138 -58 172
rect 58 138 160 172
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
rect -160 -172 -58 -138
rect 58 -172 160 -138
<< metal1 >>
rect -172 172 -46 178
rect -172 138 -160 172
rect -58 138 -46 172
rect -172 132 -46 138
rect 46 172 172 178
rect 46 138 58 172
rect 160 138 172 172
rect 46 132 172 138
rect -241 88 -195 100
rect -241 -88 -235 88
rect -201 -88 -195 88
rect -241 -100 -195 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 195 88 241 100
rect 195 -88 201 88
rect 235 -88 241 88
rect 195 -100 241 -88
rect -172 -138 -46 -132
rect -172 -172 -160 -138
rect -58 -172 -46 -138
rect -172 -178 -46 -172
rect 46 -138 172 -132
rect 46 -172 58 -138
rect 160 -172 172 -138
rect 46 -178 172 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
