magic
tech sky130A
magscale 1 2
timestamp 1729309557
<< viali >>
rect 2667 1544 2701 1578
rect 2755 1544 2789 1578
rect 942 656 976 690
rect 1066 655 1100 689
<< metal1 >>
rect 1002 2919 3043 2972
rect -25 1247 -19 1301
rect 35 1247 260 1301
rect 1002 1280 1055 2919
rect 2989 2706 3043 2919
rect 1795 2446 2007 2480
rect 1795 2103 1829 2446
rect 1658 2069 1829 2103
rect 2655 1578 2801 1584
rect 2655 1544 2667 1578
rect 2701 1544 2755 1578
rect 2789 1544 2801 1578
rect 749 1227 1055 1280
rect 1796 1507 1966 1541
rect 2655 1538 2801 1544
rect 1796 1104 1830 1507
rect 1658 1070 1830 1104
rect 930 695 988 696
rect 930 690 1112 695
rect 930 656 942 690
rect 976 689 1112 690
rect 976 656 1066 689
rect 930 655 1066 656
rect 1100 655 1112 689
rect 930 649 1112 655
<< via1 >>
rect -19 1247 35 1301
<< metal2 >>
rect -19 2972 3785 3026
rect -19 1301 35 2972
rect 3731 2677 3785 2972
rect 981 2257 990 2270
rect 828 2222 990 2257
rect 827 2135 862 2222
rect 981 2210 990 2222
rect 1050 2210 1059 2270
rect -19 1241 35 1247
<< via2 >>
rect 990 2210 1050 2270
<< metal3 >>
rect 985 2270 1055 2275
rect 985 2210 990 2270
rect 1050 2210 1437 2270
rect 985 2205 1055 2210
use differential  differential_0
timestamp 1729259257
transform 1 0 1206 0 1 2315
box -194 -1695 623 587
use ndiff  ndiff_0
timestamp 1729309557
transform 1 0 2031 0 1 2358
box -176 -1595 670 544
use nmoscs  nmoscs_0
timestamp 1729253874
transform 1 0 3043 0 1 1609
box -288 -71 976 1273
use pmoscs  pmoscs_0
timestamp 1729252742
transform 1 0 176 0 1 101
box -176 -101 836 2801
<< labels >>
flabel metal1 996 659 1020 680 0 FreeSans 800 0 0 0 vdd
port 0 nsew
flabel metal1 2709 1550 2733 1571 0 FreeSans 800 0 0 0 gnd
port 1 nsew
flabel metal1 1799 1080 1823 1101 0 FreeSans 800 0 0 0 out
port 2 nsew
flabel space 3314 2119 3338 2140 0 FreeSans 800 0 0 0 rs
port 3 nsew
flabel space 1327 2352 1351 2373 0 FreeSans 800 0 0 0 vin
port 4 nsew
flabel space 1515 2343 1539 2364 0 FreeSans 800 0 0 0 vip
port 5 nsew
<< end >>
