magic
tech sky130A
magscale 1 2
timestamp 1729309557
<< psubdiff >>
rect -176 489 -116 523
rect 610 489 670 523
rect -176 423 -142 489
rect 636 423 670 489
rect -176 -1541 -142 -1474
rect 636 -1541 670 -1474
rect -176 -1575 -116 -1541
rect 610 -1575 670 -1541
<< psubdiffcont >>
rect -116 489 610 523
rect -176 -1474 -142 423
rect 636 -1474 670 423
rect -116 -1575 610 -1541
<< poly >>
rect -30 66 0 75
rect -92 50 0 66
rect -92 16 -76 50
rect -42 16 0 50
rect -92 0 0 16
rect 494 66 524 74
rect 494 50 586 66
rect 494 16 536 50
rect 570 16 586 50
rect 494 0 586 16
rect 58 -100 436 0
rect -27 -410 0 -401
rect -92 -426 0 -410
rect -92 -460 -76 -426
rect -42 -460 0 -426
rect -92 -476 0 -460
rect 494 -410 524 -393
rect 494 -426 585 -410
rect 494 -460 535 -426
rect 569 -460 585 -426
rect 494 -476 585 -460
rect 58 -576 436 -476
rect -92 -592 0 -576
rect -92 -626 -76 -592
rect -42 -626 0 -592
rect -92 -642 0 -626
rect -29 -648 0 -642
rect 494 -592 586 -576
rect 494 -626 536 -592
rect 570 -626 586 -592
rect 494 -642 586 -626
rect 494 -664 524 -642
rect 58 -1051 436 -951
rect -92 -1067 0 -1051
rect -92 -1101 -76 -1067
rect -42 -1101 0 -1067
rect -92 -1116 0 -1101
rect 494 -1067 586 -1051
rect 494 -1101 536 -1067
rect 570 -1101 586 -1067
rect -92 -1117 -26 -1116
rect 494 -1117 586 -1101
rect 494 -1133 524 -1117
<< polycont >>
rect -76 16 -42 50
rect 536 16 570 50
rect -76 -460 -42 -426
rect 535 -460 569 -426
rect -76 -626 -42 -592
rect 536 -626 570 -592
rect -76 -1101 -42 -1067
rect 536 -1101 570 -1067
<< locali >>
rect -176 489 -116 523
rect 610 489 670 523
rect -176 423 -142 489
rect 636 423 670 489
rect -92 16 -76 50
rect -42 16 -26 50
rect 520 16 536 50
rect 570 16 586 50
rect -92 -460 -76 -426
rect -42 -460 -26 -426
rect 519 -460 535 -426
rect 569 -460 585 -426
rect -92 -626 -76 -592
rect -42 -626 -26 -592
rect 520 -626 536 -592
rect 570 -626 586 -592
rect -92 -1101 -76 -1067
rect -42 -1101 -26 -1067
rect 520 -1101 536 -1067
rect 570 -1101 586 -1067
rect -176 -1541 -142 -1474
rect 636 -1541 670 -1474
rect -176 -1575 -116 -1541
rect 610 -1575 670 -1541
<< viali >>
rect 230 489 264 523
rect -76 16 -42 50
rect 536 16 570 50
rect -76 -460 -42 -426
rect 535 -460 569 -426
rect -76 -626 -42 -592
rect 536 -626 570 -592
rect -76 -1101 -42 -1067
rect 536 -1101 570 -1067
rect 230 -1541 264 -1540
rect 230 -1575 264 -1541
<< metal1 >>
rect 211 480 221 532
rect 273 480 283 532
rect 527 443 579 449
rect -82 394 527 440
rect -82 288 -36 394
rect 75 320 201 394
rect 527 385 579 391
rect -82 88 52 288
rect 442 276 576 288
rect 211 100 221 276
rect 273 100 283 276
rect 429 100 439 276
rect 491 100 576 276
rect 442 88 576 100
rect -76 56 -42 88
rect 536 56 570 88
rect -88 50 -30 56
rect -88 16 -76 50
rect -42 16 -30 50
rect -88 10 -30 16
rect 524 50 582 56
rect 524 16 536 50
rect 570 16 582 50
rect 524 10 582 16
rect 527 -51 579 -45
rect 527 -109 579 -103
rect 530 -188 576 -109
rect -82 -200 52 -188
rect -95 -376 -85 -200
rect -33 -376 52 -200
rect 211 -376 221 -200
rect 273 -376 283 -200
rect -82 -388 52 -376
rect 442 -388 576 -188
rect -76 -420 -42 -388
rect 530 -420 576 -388
rect -88 -426 -30 -420
rect -88 -460 -76 -426
rect -42 -460 -30 -426
rect -88 -466 -30 -460
rect 523 -426 581 -420
rect 523 -460 535 -426
rect 569 -460 581 -426
rect 523 -466 581 -460
rect 530 -586 576 -466
rect -88 -592 -30 -586
rect -88 -626 -76 -592
rect -42 -626 -30 -592
rect -88 -632 -30 -626
rect 524 -592 582 -586
rect 524 -626 536 -592
rect 570 -626 582 -592
rect 524 -632 582 -626
rect -76 -664 -42 -632
rect 530 -664 576 -632
rect -82 -676 52 -664
rect -95 -852 -85 -676
rect -33 -852 52 -676
rect 211 -852 221 -676
rect 273 -852 283 -676
rect -82 -864 52 -852
rect 442 -864 576 -664
rect 530 -948 576 -864
rect 521 -1000 527 -948
rect 579 -1000 585 -948
rect -88 -1067 -30 -1061
rect -88 -1101 -76 -1067
rect -42 -1101 -30 -1067
rect -88 -1107 -30 -1101
rect 524 -1067 582 -1061
rect 524 -1101 536 -1067
rect 570 -1101 582 -1067
rect 524 -1107 582 -1101
rect -76 -1139 -42 -1107
rect 536 -1139 570 -1107
rect -82 -1339 52 -1139
rect 442 -1151 576 -1139
rect 211 -1327 221 -1151
rect 273 -1327 283 -1151
rect 429 -1327 439 -1151
rect 491 -1327 576 -1151
rect 442 -1339 576 -1327
rect -82 -1445 -36 -1339
rect 75 -1445 201 -1371
rect 527 -1442 579 -1436
rect -82 -1491 527 -1445
rect 527 -1500 579 -1494
rect 224 -1531 270 -1528
rect 211 -1583 221 -1531
rect 273 -1583 283 -1531
rect 224 -1587 270 -1583
<< via1 >>
rect 221 523 273 532
rect 221 489 230 523
rect 230 489 264 523
rect 264 489 273 523
rect 221 480 273 489
rect 527 391 579 443
rect 221 100 273 276
rect 439 100 491 276
rect 527 -103 579 -51
rect -85 -376 -33 -200
rect 221 -376 273 -200
rect -85 -852 -33 -676
rect 221 -852 273 -676
rect 527 -1000 579 -948
rect 221 -1327 273 -1151
rect 439 -1327 491 -1151
rect 527 -1494 579 -1442
rect 221 -1540 273 -1531
rect 221 -1575 230 -1540
rect 230 -1575 264 -1540
rect 264 -1575 273 -1540
rect 221 -1583 273 -1575
<< metal2 >>
rect 219 534 275 544
rect 219 468 275 478
rect -36 439 488 440
rect -82 394 488 439
rect -82 -190 -36 394
rect 442 286 488 394
rect 521 391 527 443
rect 579 391 585 443
rect 219 276 275 286
rect 219 90 275 100
rect 439 276 491 286
rect 439 90 491 100
rect 530 -51 576 391
rect 521 -103 527 -51
rect 579 -103 585 -51
rect -85 -200 -33 -190
rect -85 -386 -33 -376
rect 219 -200 275 -190
rect 219 -386 275 -376
rect -82 -666 -36 -386
rect -85 -676 -33 -666
rect -85 -862 -33 -852
rect 219 -676 275 -666
rect 219 -862 275 -852
rect -82 -1445 -36 -862
rect 527 -948 579 -942
rect 527 -1006 579 -1000
rect 219 -1151 275 -1141
rect 219 -1337 275 -1327
rect 439 -1151 491 -1141
rect 439 -1337 491 -1327
rect 442 -1445 488 -1337
rect 530 -1442 576 -1006
rect -82 -1491 488 -1445
rect 521 -1494 527 -1442
rect 579 -1494 585 -1442
rect 219 -1529 275 -1519
rect 219 -1595 275 -1585
<< via2 >>
rect 219 532 275 534
rect 219 480 221 532
rect 221 480 273 532
rect 273 480 275 532
rect 219 478 275 480
rect 219 100 221 276
rect 221 100 273 276
rect 273 100 275 276
rect 219 -376 221 -200
rect 221 -376 273 -200
rect 273 -376 275 -200
rect 219 -852 221 -676
rect 221 -852 273 -676
rect 273 -852 275 -676
rect 219 -1327 221 -1151
rect 221 -1327 273 -1151
rect 273 -1327 275 -1151
rect 219 -1531 275 -1529
rect 219 -1583 221 -1531
rect 221 -1583 273 -1531
rect 273 -1583 275 -1531
rect 219 -1585 275 -1583
<< metal3 >>
rect 209 534 285 539
rect 209 478 219 534
rect 275 478 285 534
rect 209 276 285 478
rect 209 100 219 276
rect 275 100 285 276
rect 209 95 285 100
rect 212 -195 282 95
rect 209 -200 285 -195
rect 209 -376 219 -200
rect 275 -376 285 -200
rect 209 -381 285 -376
rect 212 -671 282 -381
rect 209 -676 285 -671
rect 209 -852 219 -676
rect 275 -852 285 -676
rect 209 -857 285 -852
rect 212 -1146 282 -857
rect 209 -1151 285 -1146
rect 209 -1327 219 -1151
rect 275 -1327 285 -1151
rect 209 -1332 285 -1327
rect 210 -1524 285 -1332
rect 209 -1529 285 -1524
rect 209 -1585 219 -1529
rect 275 -1585 285 -1529
rect 209 -1590 285 -1585
use sky130_fd_pr__nfet_01v8_5MNGBB  sky130_fd_pr__nfet_01v8_5MNGBB_0
timestamp 1729238048
transform 1 0 247 0 1 -288
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGBB  sky130_fd_pr__nfet_01v8_5MNGBB_1
timestamp 1729238048
transform 1 0 247 0 1 188
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGBB  sky130_fd_pr__nfet_01v8_5MNGBB_2
timestamp 1729238048
transform 1 0 247 0 1 -1239
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_5MNGBB  sky130_fd_pr__nfet_01v8_5MNGBB_3
timestamp 1729238048
transform 1 0 247 0 1 -764
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729238506
transform 1 0 509 0 1 -1239
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729238506
transform 1 0 509 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729238506
transform 1 0 509 0 1 -288
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729238506
transform 1 0 509 0 1 -764
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1729238506
transform 1 0 -15 0 1 -1239
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1729238506
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1729238506
transform 1 0 -15 0 1 -288
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1729238506
transform 1 0 -15 0 1 -764
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_CV2X3M  XM9
timestamp 0
transform 1 0 546 0 1 -789
box 0 0 1 1
<< labels >>
flabel locali 621 501 634 509 0 FreeSans 480 0 0 0 gnd
port 0 nsew
flabel metal2 538 308 551 316 0 FreeSans 480 0 0 0 d8
port 1 nsew
flabel metal2 -67 -534 -54 -526 0 FreeSans 480 0 0 0 d9
port 2 nsew
<< end >>
