magic
tech sky130A
magscale 1 2
timestamp 1729253874
<< psubdiff >>
rect -288 1233 -228 1267
rect 916 1233 976 1267
rect -288 1211 -254 1233
rect 942 1211 976 1233
rect -288 -31 -254 -5
rect 942 -31 976 -5
rect -288 -65 -228 -31
rect 916 -65 976 -31
<< psubdiffcont >>
rect -228 1233 916 1267
rect -288 -5 -254 1211
rect 942 -5 976 1211
rect -228 -65 916 -31
<< poly >>
rect -204 1178 -112 1194
rect -204 1144 -188 1178
rect -154 1144 -112 1178
rect -204 1128 -112 1144
rect -142 1114 -112 1128
rect 800 1178 892 1194
rect 800 1144 842 1178
rect 876 1144 892 1178
rect 800 1128 892 1144
rect 800 1114 830 1128
rect 58 576 630 618
rect -142 66 -112 80
rect -204 50 -112 66
rect -204 16 -188 50
rect -154 16 -112 50
rect -204 0 -112 16
rect 800 66 830 80
rect 800 50 892 66
rect 800 16 842 50
rect 876 16 892 50
rect 800 0 892 16
<< polycont >>
rect -188 1144 -154 1178
rect 842 1144 876 1178
rect -188 16 -154 50
rect 842 16 876 50
<< locali >>
rect -288 1233 -228 1267
rect 916 1233 976 1267
rect -288 1211 -254 1233
rect 942 1211 976 1233
rect -204 1144 -188 1178
rect -154 1144 -138 1178
rect 826 1144 842 1178
rect 876 1144 892 1178
rect -204 16 -188 50
rect -154 16 -138 50
rect 826 16 842 50
rect 876 16 892 50
rect -288 -31 -254 -5
rect 942 -31 976 -5
rect -288 -65 -228 -31
rect 916 -65 976 -31
<< viali >>
rect 270 1233 304 1267
rect -188 1144 -154 1178
rect 842 1144 876 1178
rect -188 16 -154 50
rect 842 16 876 50
rect 384 -65 418 -31
<< metal1 >>
rect 258 1267 316 1273
rect 258 1233 270 1267
rect 304 1233 316 1267
rect 258 1227 316 1233
rect -200 1178 -142 1184
rect -200 1144 -188 1178
rect -154 1144 -142 1178
rect -200 1138 -142 1144
rect -188 1106 -154 1138
rect 270 1106 304 1227
rect 830 1178 888 1184
rect 830 1144 842 1178
rect 876 1144 888 1178
rect 830 1138 888 1144
rect 842 1106 876 1138
rect -194 706 52 1106
rect 264 706 310 1106
rect 378 1094 424 1106
rect 636 1094 882 1106
rect 365 718 375 1094
rect 427 718 437 1094
rect 636 718 688 1094
rect 742 718 882 1094
rect 378 706 424 718
rect 636 706 882 718
rect 12 668 46 706
rect 12 634 150 668
rect 270 618 304 706
rect 270 576 418 618
rect 384 488 418 576
rect 549 526 676 560
rect 642 488 676 526
rect -194 476 52 488
rect 265 476 310 488
rect -194 100 -54 476
rect 0 100 52 476
rect 251 100 261 476
rect 313 100 323 476
rect -194 88 52 100
rect 265 88 310 100
rect 378 88 425 488
rect 636 88 882 488
rect -188 56 -154 88
rect -200 50 -142 56
rect -200 16 -188 50
rect -154 16 -142 50
rect -200 10 -142 16
rect 384 -25 418 88
rect 842 56 876 88
rect 830 50 888 56
rect 830 16 842 50
rect 876 16 888 50
rect 830 10 888 16
rect 372 -31 430 -25
rect 372 -65 384 -31
rect 418 -65 430 -31
rect 372 -71 430 -65
<< via1 >>
rect 375 718 427 1094
rect 688 718 742 1094
rect -54 100 0 476
rect 261 100 313 476
<< metal2 >>
rect 375 1094 427 1104
rect 375 708 427 718
rect 688 1094 742 1104
rect -66 567 -57 627
rect 3 567 12 627
rect 378 620 424 708
rect 688 627 742 718
rect 264 574 424 620
rect -54 476 0 567
rect 264 486 310 574
rect 676 567 685 627
rect 745 567 754 627
rect -54 90 0 100
rect 261 476 313 486
rect 261 90 313 100
<< via2 >>
rect -57 567 3 627
rect 685 567 745 627
<< metal3 >>
rect -62 627 8 632
rect 680 627 750 632
rect -62 567 -57 627
rect 3 567 685 627
rect 745 567 750 627
rect -62 562 8 567
rect 680 562 750 567
use sky130_fd_pr__nfet_01v8_46AA6M  sky130_fd_pr__nfet_01v8_46AA6M_0
timestamp 1729217985
transform 1 0 344 0 1 597
box -344 -597 344 597
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_0
timestamp 1729217985
transform 1 0 -127 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_1
timestamp 1729217985
transform 1 0 815 0 1 906
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1729217985
transform 1 0 815 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1729217985
transform 1 0 -127 0 1 906
box -73 -226 73 226
<< labels >>
flabel locali 929 1243 943 1254 0 FreeSans 480 0 0 0 gnd
port 0 nsew
flabel metal1 -43 819 -29 830 0 FreeSans 480 0 0 0 d3
port 1 nsew
flabel metal2 705 670 719 681 0 FreeSans 480 0 0 0 d4
port 2 nsew
flabel metal2 394 654 408 665 0 FreeSans 480 0 0 0 rs
port 3 nsew
<< end >>
