magic
tech sky130A
magscale 1 2
timestamp 1729259257
<< nwell >>
rect -194 79 623 587
rect -194 58 415 79
rect 481 69 623 79
rect 418 58 623 69
rect -194 -422 623 58
rect -194 -431 -23 -422
rect -194 -456 -8 -431
rect 43 -456 623 -422
rect -194 -1695 623 -456
<< nsubdiff >>
rect -140 517 -80 551
rect 526 517 586 551
rect -140 495 -106 517
rect 552 495 586 517
rect -140 -1625 -106 -1603
rect 552 -1625 586 -1603
rect -140 -1659 -80 -1625
rect 526 -1659 586 -1625
<< nsubdiffcont >>
rect -80 517 526 551
rect -140 -1603 -106 495
rect 552 -1603 586 495
rect -80 -1659 526 -1625
<< poly >>
rect 6 69 36 80
rect -56 53 36 69
rect -56 19 -40 53
rect -6 19 36 53
rect -56 3 36 19
rect 410 69 440 85
rect 410 53 502 69
rect 410 19 452 53
rect 486 19 502 53
rect 410 3 502 19
rect 6 -431 36 -405
rect -56 -447 36 -431
rect -56 -481 -40 -447
rect -6 -481 36 -447
rect -56 -497 36 -481
rect 410 -431 440 -414
rect 410 -447 502 -431
rect 410 -481 452 -447
rect 486 -481 502 -447
rect 410 -497 502 -481
rect -56 -598 36 -582
rect -56 -632 -40 -598
rect -6 -632 36 -598
rect 94 -603 194 -497
rect 252 -603 352 -497
rect 410 -599 502 -583
rect -56 -648 36 -632
rect 6 -700 36 -648
rect 410 -633 452 -599
rect 486 -633 502 -599
rect 410 -649 502 -633
rect 410 -688 440 -649
rect -56 -1098 36 -1082
rect -56 -1132 -40 -1098
rect -6 -1132 36 -1098
rect -56 -1148 36 -1132
rect 6 -1197 36 -1148
rect 410 -1098 502 -1082
rect 410 -1132 452 -1098
rect 486 -1132 502 -1098
rect 410 -1148 502 -1132
rect 410 -1187 440 -1148
<< polycont >>
rect -40 19 -6 53
rect 452 19 486 53
rect -40 -481 -6 -447
rect 452 -481 486 -447
rect -40 -632 -6 -598
rect 452 -633 486 -599
rect -40 -1132 -6 -1098
rect 452 -1132 486 -1098
<< locali >>
rect -140 517 -80 551
rect 526 517 586 551
rect -140 495 -106 517
rect 552 495 586 517
rect -56 19 -40 53
rect -6 19 10 53
rect 436 19 452 53
rect 486 19 502 53
rect -56 -481 -40 -447
rect -6 -481 10 -447
rect 436 -481 452 -447
rect 486 -481 502 -447
rect -56 -632 -40 -598
rect -6 -632 10 -598
rect 436 -633 452 -599
rect 486 -633 502 -599
rect -56 -1132 -40 -1098
rect -6 -1132 10 -1098
rect 436 -1132 452 -1098
rect 486 -1132 502 -1098
rect -140 -1625 -106 -1603
rect 552 -1625 586 -1603
rect -140 -1659 -80 -1625
rect 526 -1659 586 -1625
<< viali >>
rect -40 19 -6 53
rect 452 19 486 53
rect -40 -481 -6 -447
rect 452 -481 486 -447
rect -40 -632 -6 -598
rect 452 -633 486 -599
rect -40 -1132 -6 -1098
rect 452 -1132 486 -1098
rect 197 -1388 249 -1212
<< metal1 >>
rect 443 464 495 470
rect -46 415 443 461
rect -46 300 0 415
rect 443 406 495 412
rect -46 100 88 300
rect 358 288 492 300
rect 187 112 197 288
rect 249 112 259 288
rect 345 112 355 288
rect 407 112 492 288
rect 358 100 492 112
rect -40 59 -6 100
rect -52 53 6 59
rect -52 19 -40 53
rect -6 19 6 53
rect -52 13 6 19
rect 100 10 110 62
rect 178 10 188 62
rect 452 59 486 100
rect 440 53 498 59
rect 268 -19 336 53
rect 440 19 452 53
rect 486 19 498 53
rect 440 13 498 19
rect 110 -81 336 -19
rect 110 -132 178 -81
rect 443 -110 495 -104
rect 258 -162 268 -110
rect 336 -162 346 -110
rect 443 -168 495 -162
rect 446 -200 492 -168
rect -46 -212 88 -200
rect -59 -388 -49 -212
rect 3 -388 88 -212
rect 187 -388 197 -212
rect 249 -388 259 -212
rect -46 -400 88 -388
rect 358 -400 492 -200
rect -40 -441 -6 -400
rect 446 -441 492 -400
rect -52 -447 6 -441
rect -52 -481 -40 -447
rect -6 -481 6 -447
rect -52 -487 6 -481
rect 440 -447 498 -441
rect 440 -481 452 -447
rect 486 -481 498 -447
rect 440 -487 498 -481
rect -52 -598 6 -592
rect 446 -593 492 -487
rect -52 -632 -40 -598
rect -6 -632 6 -598
rect -52 -638 6 -632
rect 440 -599 498 -593
rect 440 -633 452 -599
rect 486 -633 498 -599
rect -40 -700 -6 -638
rect 440 -639 498 -633
rect 446 -700 492 -639
rect -46 -712 88 -700
rect -59 -888 -49 -712
rect 3 -888 88 -712
rect 187 -888 197 -712
rect 249 -888 259 -712
rect -46 -900 88 -888
rect 358 -900 492 -700
rect 446 -938 492 -900
rect 100 -990 110 -938
rect 178 -990 188 -938
rect 268 -1019 336 -981
rect 437 -990 443 -938
rect 495 -990 501 -938
rect 110 -1081 336 -1019
rect -52 -1098 6 -1092
rect -52 -1132 -40 -1098
rect -6 -1132 6 -1098
rect 110 -1127 178 -1081
rect 440 -1098 498 -1092
rect -52 -1138 6 -1132
rect -40 -1200 -6 -1138
rect 258 -1162 268 -1110
rect 336 -1162 346 -1110
rect 440 -1132 452 -1098
rect 486 -1132 498 -1098
rect 440 -1138 498 -1132
rect 452 -1200 486 -1138
rect -46 -1400 88 -1200
rect 191 -1212 255 -1200
rect 358 -1212 492 -1200
rect 187 -1388 197 -1212
rect 249 -1388 259 -1212
rect 345 -1388 355 -1212
rect 407 -1388 492 -1212
rect 191 -1400 255 -1388
rect 358 -1400 492 -1388
rect -46 -1515 0 -1400
rect 443 -1512 495 -1506
rect -46 -1561 443 -1515
rect 443 -1570 495 -1564
<< via1 >>
rect 443 412 495 464
rect 197 112 249 288
rect 355 112 407 288
rect 110 10 178 62
rect 268 -162 336 -110
rect 443 -162 495 -110
rect -49 -388 3 -212
rect 197 -388 249 -212
rect -49 -888 3 -712
rect 197 -888 249 -712
rect 110 -990 178 -938
rect 443 -990 495 -938
rect 268 -1162 336 -1110
rect 197 -1388 249 -1212
rect 355 -1388 407 -1212
rect 443 -1564 495 -1512
<< metal2 >>
rect -46 415 404 461
rect -46 -202 0 415
rect 358 298 404 415
rect 437 412 443 464
rect 495 412 501 464
rect 195 288 251 298
rect 195 102 251 112
rect 355 288 407 298
rect 355 102 407 112
rect 110 62 178 72
rect 110 3 178 10
rect 110 -103 336 3
rect 268 -110 336 -103
rect 446 -110 492 412
rect 437 -162 443 -110
rect 495 -162 501 -110
rect 268 -172 336 -162
rect -49 -212 3 -202
rect -49 -398 3 -388
rect 195 -212 251 -202
rect 195 -398 251 -388
rect -46 -702 0 -398
rect -49 -712 3 -702
rect -49 -898 3 -888
rect 195 -712 251 -702
rect 195 -898 251 -888
rect -46 -1515 0 -898
rect 110 -938 178 -928
rect 110 -997 178 -990
rect 443 -938 495 -932
rect 443 -996 495 -990
rect 110 -1103 336 -997
rect 268 -1110 336 -1103
rect 268 -1172 336 -1162
rect 195 -1212 251 -1202
rect 195 -1398 251 -1388
rect 355 -1212 407 -1202
rect 355 -1398 407 -1388
rect 358 -1515 404 -1398
rect 446 -1512 492 -996
rect -46 -1561 404 -1515
rect 437 -1564 443 -1512
rect 495 -1564 501 -1512
<< via2 >>
rect 195 112 197 288
rect 197 112 249 288
rect 249 112 251 288
rect 195 -388 197 -212
rect 197 -388 249 -212
rect 249 -388 251 -212
rect 195 -888 197 -712
rect 197 -888 249 -712
rect 249 -888 251 -712
rect 195 -1388 197 -1212
rect 197 -1388 249 -1212
rect 249 -1388 251 -1212
<< metal3 >>
rect 185 288 261 293
rect 185 112 195 288
rect 251 112 261 288
rect 185 -212 261 112
rect 185 -388 195 -212
rect 251 -388 261 -212
rect 185 -712 261 -388
rect 185 -888 195 -712
rect 251 -888 261 -712
rect 185 -1212 261 -888
rect 185 -1388 195 -1212
rect 251 -1388 261 -1212
rect 185 -1393 261 -1388
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729231080
transform 1 0 21 0 1 -800
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729231080
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729231080
transform 1 0 425 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729231080
transform 1 0 425 0 1 -800
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729231080
transform 1 0 425 0 1 -1300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729231080
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729231080
transform 1 0 21 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729231080
transform 1 0 21 0 1 -1300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_0
timestamp 1729228836
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_1
timestamp 1729228836
transform 1 0 223 0 1 -300
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_2
timestamp 1729228836
transform 1 0 223 0 1 -800
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXXLL  sky130_fd_pr__pfet_01v8_VQXXLL_3
timestamp 1729228836
transform 1 0 223 0 1 -1300
box -223 -200 223 200
<< labels >>
flabel metal3 205 -526 217 -520 0 FreeSans 480 0 0 0 s
port 1 nsew
flabel metal2 134 -10 146 -4 0 FreeSans 480 0 0 0 vin
port 2 nsew
flabel metal1 277 35 289 41 0 FreeSans 480 0 0 0 vip
port 3 nsew
flabel metal2 375 354 387 360 0 FreeSans 480 0 0 0 d7
port 4 nsew
flabel metal2 470 -62 482 -56 0 FreeSans 480 0 0 0 d6
port 5 nsew
flabel locali 544 529 556 535 0 FreeSans 480 0 0 0 vdd
port 0 nsew
<< end >>
